`timescale 1ns / 1ps

module ffd_tb;


//declaration of signals
parameter W = 5;
reg clk; //system clock
reg rst; //system reset
reg enable; //load signal
reg [W-1:0] D; //input signal
wire [W-1:0] Q; //output signal

//Instantiation of the D flip flop
d_ff_en	#(.W(W)) dut 
(
	.clk(clk), 			//system clock
	.rst(rst), 			//system reset
	.enable(enable),	//load signal
	.D(D), 				//input signal
	.Q(Q)				//output signal
);

//Generation of the clock
initial begin
	clk = 0;
	forever #5 clk = ~clk;
end

//Stimulus specification

initial
begin
	#100
	rst = 1;
	enable = 0;
	D = 5'b00000;
	#10
	rst = 0;
	enable = 1;

	#10
	D = 5'b11001;

	#10
	enable = 0;

	#10
	D = 5'b11111;

	#30
	enable = 1;

	#20
	rst = 1;

	#30 $stop;
end

integer f,i;

initial
begin
f=$fopen("output.txt","w");
$timeformat(-9,1,"ns",12);
$display(" 	Time 	clk 	rst	 EN	 D 	Q");
$monitor("%t %b %b %b %b %b", $realtime,clk,rst,enable,D,Q);
for(i=0; i<44;i=i+1)
begin
@(clk)
$fwrite(f,"%t %b %b %b %b %b\n", $realtime,clk,rst,enable,D,Q);
end
$fclose(f);

end

endmodule
